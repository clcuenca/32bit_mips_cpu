library verilog;
use verilog.vl_types.all;
entity mips_32_vlg_vec_tst is
end mips_32_vlg_vec_tst;
