library verilog;
use verilog.vl_types.all;
entity data_memory_4kb is
    port(
        clock           : in     vl_logic;
        memread         : in     vl_logic;
        memwrite        : in     vl_logic;
        address         : in     vl_logic_vector(31 downto 0);
        write_data      : in     vl_logic_vector(31 downto 0);
        read_data       : out    vl_logic_vector(31 downto 0)
    );
end data_memory_4kb;
