library verilog;
use verilog.vl_types.all;
entity mips_32 is
    port(
        clock           : in     vl_logic
    );
end mips_32;
